module register(q, d, wrenable, clk);
  input d;
  input wrenable;
  input clk;
  output reg q;
  always @(posedge clk) begin
    if(wrenable) begin
      q = d;
    end
  end
endmodule

module register32(q, d, wrenable, clk);
  parameter busWidth = 32;
  input[busWidth - 1:0] d;
  input wrenable;
  input clk;
  output reg[busWidth - 1:0] q;
  always @(posedge clk) begin
    if(wrenable) begin
      q = d;
    end
  end
endmodule

module register32Zero(q, d, wrenable, clk);
  parameter busWidth = 32;
  input[busWidth - 1:0] d;
  input wrenable;
  input clk;
  output reg[busWidth - 1:0] q;
  always @(posedge clk) begin
      //save gates by not checking wrenable
      q = 0;
  end
endmodule

module mux32to1by1(out, address, inputs);
  input[31:0] inputs;
  input[4:0] address;
  output out;

  assign out = inputs[address];

endmodule

module mux32to1by32(out, address, input0, input1, input2, input3, input4, input5, input6, input7, input8, input9, input10, input11, input12, input13, input14, input15, input16, input17, input18, input19, input20, input21, input22, input23, input24, input25, input26, input27, input28, input29, input30, input31);
  input[31:0] input0, input1, input2, input3, input4, input5, input6, input7, input8, input9, input10, input11, input12, input13, input14, input15, input16, input17, input18, input19, input20, input21, input22, input23, input24, input25, input26, input27, input28, input29, input30, input31;
  input[4:0] address;
  output[31:0] out;
  wire[31:0] mux[31:0]; // Creates a 2d Array of wires
  assign mux[0] = input0; // Connects the sources of the array
  assign mux[1] = input1;
  assign mux[2] = input2;
  assign mux[3] = input3;
  assign mux[4] = input4;
  assign mux[5] = input5;
  assign mux[6] = input6;
  assign mux[7] = input7;
  assign mux[8] = input8;
  assign mux[9] = input9;
  assign mux[10] = input10;
  assign mux[11] = input11;
  assign mux[12] = input12;
  assign mux[13] = input13;
  assign mux[14] = input14;
  assign mux[15] = input15;
  assign mux[16] = input16;
  assign mux[17] = input17;
  assign mux[18] = input18;
  assign mux[19] = input19;
  assign mux[20] = input20;
  assign mux[21] = input21;
  assign mux[22] = input22;
  assign mux[23] = input23;
  assign mux[24] = input24;
  assign mux[25] = input25;
  assign mux[26] = input26;
  assign mux[27] = input27;
  assign mux[28] = input28;
  assign mux[29] = input29;
  assign mux[30] = input30;
  assign mux[31] = input31;

  assign out = mux[address]; // Connects the output of the array
endmodule

module decoder1to32(out, enable, address);
  output[31:0] out;
  input enable;
  input[4:0] address;
  // The "<<" operator shifts the 1 or 0 enable left by the value of the address.
  // The address can be from 0-31 and and if the enable is set to 1,
  // the decoder will therefor set the output to a 32 bit bus
  // with 1 at the bit numbered by the address with the rest of the bits 0.
  assign out = enable<<address; 
endmodule

module regfile(ReadData1, // Contents of first register read
 ReadData2, // Contents of second register read
 WriteData, // Contents to write to register
 ReadRegister1, // Address of first register to read 
 ReadRegister2, // Address of second register to read
 WriteRegister, // Address of register to write
 RegWrite, // Enable writing of register when High
 Clk); // Clock (Positive Edge Triggered)
  output[31:0] ReadData1, ReadData2;
  input[31:0] WriteData;
  input[4:0] ReadRegister1, ReadRegister2, WriteRegister;
  input RegWrite, Clk;

  wire[31:0] regWriteIndex;
  wire[31:0] regOuts[31:0];
  decoder1to32 decoder(regWriteIndex, RegWrite, WriteRegister);
  register32Zero reg0(regOuts[0], WriteData, regWriteIndex[0], Clk);
  generate
    genvar i;
    for (i = 1; i < 32; i = i + 1) begin
      register32 reg1(regOuts[i], WriteData, regWriteIndex[i], Clk);
    end
  endgenerate
  mux32to1by32 mux1(ReadData1, ReadRegister1, regOuts[0], regOuts[1], regOuts[2], regOuts[3], regOuts[4], regOuts[5], regOuts[6], regOuts[7], regOuts[8], regOuts[9], regOuts[10], regOuts[11], regOuts[12], regOuts[13], regOuts[14], regOuts[15], regOuts[16], regOuts[17], regOuts[18], regOuts[19], regOuts[20], regOuts[21], regOuts[22], regOuts[23], regOuts[24], regOuts[25], regOuts[26], regOuts[27], regOuts[28], regOuts[29], regOuts[30], regOuts[31]);
  mux32to1by32 mux2(ReadData2, ReadRegister2, regOuts[0], regOuts[1], regOuts[2], regOuts[3], regOuts[4], regOuts[5], regOuts[6], regOuts[7], regOuts[8], regOuts[9], regOuts[10], regOuts[11], regOuts[12], regOuts[13], regOuts[14], regOuts[15], regOuts[16], regOuts[17], regOuts[18], regOuts[19], regOuts[20], regOuts[21], regOuts[22], regOuts[23], regOuts[24], regOuts[25], regOuts[26], regOuts[27], regOuts[28], regOuts[29], regOuts[30], regOuts[31]);

endmodule

// Validates your hw4testbench by connecting it to various functional 
// or broken register files and verifying that it correctly identifies 
module regfiletestbenchharness;
wire[31:0]  ReadData1;
wire[31:0]  ReadData2;
wire[31:0]  WriteData;
wire[4:0] ReadRegister1;
wire[4:0] ReadRegister2;
wire[4:0] WriteRegister;
wire    RegWrite;
wire    Clk;
reg   begintest;

// The register file being tested.  DUT = Device Under Test
regfile DUT(ReadData1, ReadData2, WriteData, ReadRegister1, ReadRegister2, WriteRegister, RegWrite, Clk);

// The test harness to test the DUT
hw4testbench tester(begintest, endtest, dutpassed, ReadData1,ReadData2,WriteData, ReadRegister1, ReadRegister2, WriteRegister, RegWrite, Clk);


initial begin
begintest=0;
#10;
begintest=1;
#1000;
end

always @(posedge endtest) begin
$display(dutpassed);
end

endmodule

// This is your
// It generates the signals to drive a registerfile and passes it back up one layer to the harness
//  ((This lets us plug in various working / broken registerfiles to test
// When begintest is asserted, begin testing the register file.
// When your test is conclusive, set dutpassed as appropriate and then raise endtest.
module regfiletestbench(begintest, endtest, dutpassed,
        ReadData1,ReadData2,WriteData, ReadRegister1, ReadRegister2,WriteRegister,RegWrite, Clk);
output reg endtest;
output reg dutpassed;
input    begintest;

input[31:0]   ReadData1;
input[31:0]   ReadData2;
output reg[31:0]  WriteData;
output reg[4:0]   ReadRegister1;
output reg[4:0]   ReadRegister2;
output reg[4:0]   WriteRegister;
output reg    RegWrite;
output reg    Clk;

initial begin
WriteData=0;
ReadRegister1=0;
ReadRegister2=0;
WriteRegister=0;
RegWrite=0;
Clk=0;
end

always @(posedge begintest) begin
endtest = 0;
dutpassed = 1;
#10

// Test Case 1: Write 42 to register 2, verify with Read Ports 1 and 2
// This will pass because the example register file is hardwired to always return 42.
WriteRegister = 2;
WriteData = 42;
RegWrite = 1;
ReadRegister1 = 2;
ReadRegister2 = 2;
#5 Clk=1; #5 Clk=0; // Generate Clock Edge
if(ReadData1 != 42 || ReadData2!= 42) begin
  dutpassed = 0;
  $display("Test Case 1 Failed");
  end

// Test Case 2: Write 15 to register 2, verify with Read Ports 1 and 2
// This will fail with the example register file, but should pass with yours.
WriteRegister = 2;
WriteData = 15;
RegWrite = 1;
ReadRegister1 = 2;
ReadRegister2 = 2;
#5 Clk=1; #5 Clk=0;
if(ReadData1 != 15 || ReadData2!= 15) begin
  dutpassed = 0;  // On Failure, set to false.
  $display("Test Case 2 Failed");
  end


// Test Case 3: Test WriteEnable blocks writes when off
// Write 16 to register 2, verify with Read Ports 1 and 2
WriteRegister = 2;
WriteData = 16;
RegWrite = 0;
ReadRegister1 = 2;
ReadRegister2 = 2;
#5 Clk=1; #5 Clk=0;
if(ReadData1 == 16 || ReadData2 == 16) begin
  dutpassed = 0;  // On Failure, set to false.
  $display("Test Case 3 Failed, WriteEnable does not control writing.");
  end

// Test Case 4: Test Decoder specifies writing to a single register
// Write 18 to register 2, verify with Read Ports 1 and 2
WriteRegister = 2;
WriteData = 18;
RegWrite = 1;
ReadRegister1 = 4;
ReadRegister2 = 4;
#5 Clk=1; #5 Clk=0;
if(ReadData1 == 18 || ReadData2 == 18) begin
  dutpassed = 0;  // On Failure, set to false.
  $display("Test Case 4 Failed, Non-targeted register written to.");
  end

// Test Case 5: Test registerZero is not writable
// Write 4 to register 0, verify with Read Ports 1 and 2
WriteRegister = 0;
WriteData = 4;
RegWrite = 1;
ReadRegister1 = 0;
ReadRegister2 = 0;
#5 Clk=1; #5 Clk=0;
if(ReadData1 == 4 || ReadData2 == 4) begin
  dutpassed = 0;  // On Failure, set to false.
  $display("Test Case 5 Failed, Register 0 is writable.");
  end

// Test Case 6: Test registerZero contains value zero
// Read register zero
WriteRegister = 0;
WriteData = 4;
RegWrite = 1;
ReadRegister1 = 0;
ReadRegister2 = 0;
#5 Clk=1; #5 Clk=0;
if(ReadData1 != 0 || ReadData2 != 0) begin
  dutpassed = 0;  // On Failure, set to false.
  $display("Test Case 6 Failed, Register 0 does not contain zero");
  end

// Test Case 7: Test Port 2 reads correct port
// Write 12 to register 17, verify register 17 equals 12 with Port 1
// verify Port 2 reads 12 while assigned to read register 0
WriteRegister = 17;
WriteData = 12;
RegWrite = 1;
ReadRegister1 = 17;
ReadRegister2 = 0;
#5 Clk=1; #5 Clk=0;
if(ReadData1 != 12 || ReadData2 == 12) begin
  dutpassed = 0;  // On Failure, set to false.
  $display("Test Case 7 Failed, Port 2 read incorrect register.");
  end

//We're done!  Wait a moment and signal completion.
#5
endtest = 1;
end

endmodule